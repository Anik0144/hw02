magic
tech sky130A
magscale 1 2
timestamp 1680143486
<< error_p >>
rect -77 831 -19 837
rect 115 831 173 837
rect -77 797 -65 831
rect 115 797 127 831
rect -77 791 -19 797
rect 115 791 173 797
<< nwell >>
rect -161 812 257 850
rect -257 -812 257 812
rect -257 -850 161 -812
rect -190 -853 100 -850
<< pmos >>
rect -159 -750 -129 750
rect -63 -750 -33 750
rect 33 -750 63 750
rect 129 -750 159 750
<< pdiff >>
rect -221 738 -159 750
rect -221 -738 -209 738
rect -175 -738 -159 738
rect -221 -750 -159 -738
rect -129 738 -63 750
rect -129 -738 -113 738
rect -79 -738 -63 738
rect -129 -750 -63 -738
rect -33 738 33 750
rect -33 -738 -17 738
rect 17 -738 33 738
rect -33 -750 33 -738
rect 63 738 129 750
rect 63 -738 79 738
rect 113 -738 129 738
rect 63 -750 129 -738
rect 159 738 221 750
rect 159 -738 175 738
rect 209 -738 221 738
rect 159 -750 221 -738
<< pdiffc >>
rect -209 -738 -175 738
rect -113 -738 -79 738
rect -17 -738 17 738
rect 79 -738 113 738
rect 175 -738 209 738
<< poly >>
rect -81 831 -15 847
rect -81 797 -65 831
rect -31 797 -15 831
rect -81 781 -15 797
rect 111 831 177 847
rect 111 797 127 831
rect 161 797 177 831
rect 111 781 177 797
rect -159 750 -129 776
rect -63 750 -33 781
rect 33 750 63 776
rect 129 750 159 781
rect -159 -777 -129 -750
rect -63 -776 -33 -750
rect 33 -777 63 -750
rect 129 -776 159 -750
<< polycont >>
rect -65 797 -31 831
rect 127 797 161 831
<< locali >>
rect -81 797 -65 831
rect -31 797 -15 831
rect 111 797 127 831
rect 161 797 177 831
rect -209 738 -175 754
rect -209 -754 -175 -738
rect -113 738 -79 754
rect -113 -754 -79 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 79 738 113 754
rect 79 -754 113 -738
rect 175 738 209 754
rect 175 -754 209 -738
<< viali >>
rect -65 797 -31 831
rect 127 797 161 831
rect -209 -738 -175 738
rect -113 -738 -79 738
rect -17 -738 17 738
rect 79 -738 113 738
rect 175 -738 209 738
<< metal1 >>
rect -77 831 -19 837
rect -77 797 -65 831
rect -31 797 -19 831
rect -77 791 -19 797
rect 115 831 173 837
rect 115 797 127 831
rect 161 797 173 831
rect 115 791 173 797
rect -215 738 -169 750
rect -215 -738 -209 738
rect -175 -738 -169 738
rect -215 -750 -169 -738
rect -119 738 -73 750
rect -119 -738 -113 738
rect -79 -738 -73 738
rect -119 -750 -73 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 73 738 119 750
rect 73 -738 79 738
rect 113 -738 119 738
rect 73 -750 119 -738
rect 169 738 215 750
rect 169 -738 175 738
rect 209 -738 215 738
rect 169 -750 215 -738
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.5 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
